-- Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 16.0.0 Build 211 04/27/2016 SJ Lite Edition
-- Created on Thu Dec 01 17:14:33 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY FinalProject IS
    PORT (
        reset : IN STD_LOGIC := '0';
		  r : IN STD_LOGIC := '0';
		  clockState : IN STD_LOGIC;
        clock : IN STD_LOGIC;
		  Change : IN STD_LOGIC := '0';
        M500 : IN STD_LOGIC := '0';
        M1000 : IN STD_LOGIC := '0';
        T : OUT STD_LOGIC;
        Ca : OUT STD_LOGIC;
		  Display : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		  SEGMENTS : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		  Position: out std_logic
    );
	 
END FinalProject;

ARCHITECTURE BEHAVIOR OF FinalProject IS
    TYPE type_fstate IS (State0,State1500,State2000,State3000,State2500,State500,State1000);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
	 SIGNAL Transistor1, Transistor2, Transistor3, Transistor4: STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
	 SIGNAL Count : integer range 0 to 100000;
	 SIGNAL Selection : STD_LOGIC_VECTOR(1 DOWNTO 0) :="00";
	 SIGNAL toShow : STD_LOGIC_VECTOR(3 DOWNTO 0) :="0000";
	 
BEGIN

    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;
	 
	 
	 COUNTING_CLK_STATE: PROCESS(clockState)
		BEGIN
			IF RISING_EDGE(clockState) THEN
				IF Count < 100000 THEN 
				
					Count <= Count+1;
				ELSE
					Selection <= Selection+1;
					Count <= 0;
				END IF;
			END IF;
			
		END PROCESS;
	 
	 
	 	SHOW_SEGMENTS: PROCESS(Selection)
		BEGIN
			CASE Selection is
						WHEN "00"=> 
							toShow <= "1110";
							
						WHEN "01" => 
							toShow <= "1101";
							
						WHEN "10"=> 
							toShow <= "1011";
							
						WHEN "11" => 
							toShow <= "0111";
						
					   WHEN OTHERS => 
							toshow <= "1111";
							
			END CASE;
	 
	 CASE toShow is 
						
						WHEN "1110" =>
							Segments <= Transistor1;
							
						WHEN "1101" =>
							Segments <= Transistor2;
							
						WHEN "1011" =>
							Segments <= Transistor3;
							
						WHEN "0111" =>
							Segments <= Transistor4;
							
						WHEN OTHERS => 
							Segments <= "1111111";	
			END CASE;
			
		END PROCESS;
		
		Display <= toShow;
	 

    PROCESS (fstate,reset,M500,M1000)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= State0;
            T <= '0';
            Ca <= '0';
        ELSE
            T <= '0';
            Ca <= '0';
            CASE fstate IS
                WHEN State0 =>
					 
					      Transistor4 <= "0000001"; 
							Transistor3 <= "0000001"; 
							Transistor2 <= "0000001"; 
							Transistor1 <= "0000001";
							
						  T <= '0';

                    Ca <= '0';
					 
                    IF (((M500 = '0') AND (M1000 = '1'))) THEN
                        reg_fstate <= State1000;
                    ELSIF (((M500 = '1') AND (M1000 = '0'))) THEN
                        reg_fstate <= State500;
                    ELSIF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State0;
                    END IF;

                    
                WHEN State1500 =>
					 
					 
					     Transistor4 <= "0000001";
						  Transistor3 <= "0000001";
						  Transistor2 <= "0100100"; --5
						  Transistor1 <= "1001111"; --1
						  
						  T <= '0';

                    Ca <= '0';
					 
                    IF (((M500 = '0') AND (M1000 = '1'))) THEN
                        reg_fstate <= State2500;
                    ELSIF (((M500 = '1') AND (M1000 = '0'))) THEN
                        reg_fstate <= State2000;
                    ELSIF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State1500;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State1500;
                    END IF;

                   
                WHEN State2000 =>
					 
					     Transistor4 <= "0000001";
						  Transistor3 <= "0000001";
						  Transistor2 <= "0000001";
						  Transistor1 <= "0010010";
					 
					 
					     T <= '0';

                    Ca <= '0';
					 
                    IF (((M500 = '0') AND (M1000 = '1'))) THEN
                        reg_fstate <= State3000;
                    ELSIF (((M500 = '1') AND (M1000 = '0'))) THEN
                        reg_fstate <= State2500;
                    ELSIF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State2000;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State2000;
                    END IF;


                WHEN State3000 =>
					 
					     T <= '1';

                    Ca <= '1';
					  
					     Transistor4 <= "0000001";
						  Transistor3 <= "0000001";
						  Transistor2 <= "0000001";
						  Transistor1 <= "0000110";
					 
                    IF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State500;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State3000;
                    END IF;

                    
                WHEN State2500 =>
					 
					     T <= '1';

                    Ca <= '0';
					 
					     Transistor4 <= "0000001";
						  Transistor3 <= "0000001";
						  Transistor2 <= "0100100";
						  Transistor1 <= "0010010";
					 
                    IF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State0;
                    ELSIF (((M500 = '1') AND (M1000 = '0'))) THEN
                        reg_fstate <= State3000;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State2500;
                    END IF;

                    
                WHEN State500 =>
					 
					     T <= '0';

                    Ca <= '0';
					 
					     Transistor4 <= "0000001";
						  Transistor3 <= "0000001";
						  Transistor2 <= "0100100";
						  Transistor1 <= "0000001";
					 
                    IF (((M500 = '0') AND (M1000 = '1'))) THEN
                        reg_fstate <= State1500;
                    ELSIF (((M500 = '1') AND (M1000 = '0'))) THEN
                        reg_fstate <= State1000;
                    ELSIF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State500;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State500;
                    END IF;

                    
						  
                WHEN State1000 =>
					 
					     T <= '0';

                    Ca <= '0';
					 
					 
					     Transistor4 <= "0000001";
						  Transistor3 <= "0000001";
						  Transistor2 <= "0000001";
						  Transistor1 <= "1001111";
					 
					 
                    IF (((M500 = '1') AND (M1000 = '0'))) THEN
                        reg_fstate <= State1500;
                    ELSIF (((M500 = '0') AND (M1000 = '1'))) THEN
                        reg_fstate <= State2000;
                    ELSIF (((M500 = '0') AND (M1000 = '0'))) THEN
                        reg_fstate <= State1000;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State1000;
                    END IF;

                    
                WHEN OTHERS => 
					 
					     T <= 'X';
                    Ca <= 'X';
					 
					      Transistor4 <= "0000001"; 
							Transistor3 <= "0000001"; 
							Transistor2 <= "0000001"; 
							Transistor1 <= "0000001";
					 
                    
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
